library IEEE;
use IEEE.std_logic_1164.all;
library gate_lib;

entity mux_hmwk1 is
  port(a       : in std_logic;
       b       : in std_logic;
       sel     : in std_logic;
       y : out std_logic);
end mux_hmwk1;

architecture structural of mux_hmwk1 is
  
  --component declarations
  component and2 is
    generic(Tp : time := 2 ns);
    port(in1  : in std_logic;
         in2  : in std_logic;
         out1 : out std_logic);
  end component;
  
  component or2 is
    generic(Tp : time := 2 ns);
    port(in1  : in std_logic;
         in2  : in std_logic;
         out1 : out std_logic);
  end component;
  
  component inv is
    generic(Tp : time := 1 ns);
    port(in1  : in std_logic;
         out1 : out std_logic);
  end component;

  for all : and2 use entity gate_lib.and2(simple);
  for all : or2 use entity gate_lib.or2(simple);
  for all : inv use entity gate_lib.inv(simple);

  --signal statements
  signal sig_1,  sig_2,  sig_3 : std_logic;
  
  begin
    --structural descriptions
    NOT_1 : inv generic map(Tp => 1 ns)
                port map(in1 => sel,
                        out1 => sig_1);
                        
    AND_1 : and2 generic map(Tp => 2 ns)
                 port map(in1 => a, in2 => sig_1,
                        out1 => sig_2);                        
                        
    AND_2 : and2 generic map(Tp => 2 ns)
                 port map(in1 => b, in2 => sel,
                        out1 => sig_3);                     
                        
    OR_1 : or2 generic map(Tp => 2 ns)
               port map(in1 => sig_2, in2 => sig_3,
                        out1 => y);                                              
end structural;